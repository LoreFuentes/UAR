Library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;	 

entity Deserializer is
	generic(busWidth : integer := 10);
	port(
		RST : in std_logic;
		CLK : in std_logic; 
		BIN : in std_logic;
		SHF : in std_logic;
		DOUT : out std_logic_vector(busWidth-1 downto 0)
		);
end Deserializer;	   

architecture Behavioral of Deserializer is 
signal Qp,Qn : std_logic_vector(busWidth-1 downto 0);
begin

	combinatorial : process (Qp,SHF,BIN)
	begin 
		if SHF = '1' then 
			Qn <= Qp(busWidth-2 downto 0) & BIN;
		else 
			Qn <= Qp;  
		end if;
		
	DOUT <= Qp;
	end process combinatorial ;
	
	Sequential : process(RST,CLK)
	begin
		if RST = '0' then 
			Qp <= (others => '0');
		elsif  CLK' event and CLK = '1' then
			Qp <= Qn;
		end if;
	end process Sequential;
	
end Behavioral;

